-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 184 04/29/2009 Service Pack 1 SJ Web Edition
-- Created on Sat Nov 16 19:59:52 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY RCRstate IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        nrxf : IN STD_LOGIC := '0';
        ntxe : IN STD_LOGIC := '0';
        nrd : OUT STD_LOGIC;
        wr : OUT STD_LOGIC;
        din : IN STD_LOGIC_VECTOR(7 downto 0);
        dout: OUT STD_LOGIC_VECTOR(7 downto 0)
    );
END RCRstate;

ARCHITECTURE BEHAVIOR OF RCRstate IS
    TYPE type_fstate IS (wait_nrxf_low,wait_ntxe_low,set_wr_high,set_nrd_low,latch_data_from_host,send_data_host);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL o : std_logic_vector(4 downto 0);
    SIGNAL input : std_logic_vector(13 downto 0);
    SIGNAL p : std_logic_vector(5 downto 0);
    SIGNAL a_in : std_logic_vector(8 downto 0);
    SIGNAL b_out : std_logic_vector(4 downto 0);
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= wait_nrxf_low;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (clock)
    BEGIN
        nrd <= '0';
        wr <= '0';
        IF clock'event and clock='1' THEN
        CASE fstate IS
            WHEN wait_nrxf_low =>
                IF ((nrxf = '1')) THEN
                    reg_fstate <= wait_nrxf_low;
                ELSIF (NOT((nrxf = '1'))) THEN
                    reg_fstate <= set_nrd_low;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= wait_nrxf_low;
                END IF;

                nrd <= '1';

                wr <= '0';
            WHEN set_nrd_low =>
                reg_fstate <= latch_data_from_host;

                nrd <= '0';

                wr <= '0';
            WHEN latch_data_from_host =>
                reg_fstate <= wait_ntxe_low;

                nrd <= '0';

                wr <= '0';
                a_in(7 downto 0) <= din(7 downto 0);
            WHEN wait_ntxe_low =>
                IF ((ntxe = '1')) THEN
                    reg_fstate <= wait_ntxe_low;
                ELSIF (NOT((ntxe = '1'))) THEN
                    reg_fstate <= set_wr_high;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= wait_ntxe_low;
                END IF;

                nrd <= '1';

                wr <= '0';
            WHEN set_wr_high =>
                reg_fstate <= send_data_host;

                nrd <= '1';

                wr <= '1';
            WHEN send_data_host =>
                reg_fstate <= wait_nrxf_low;

                nrd <= '1';

                wr <= '1';
                dout(4 downto 0) <= o(4 downto 0);
                dout(7 downto 5) <= "000";
            WHEN OTHERS => 
                nrd <= '1';
                wr <= '1';
				dout <= "ZZZZZZZZ";
                reg_fstate <= wait_nrxf_low;
        END CASE;
        END IF;
    END PROCESS;
    
    process(clock)
	variable d: std_logic_vector(5 downto 0);
	variable c: std_logic_vector(4 downto 0);
	begin
		p <= "110101";
		c := "00000";
		input <= a_in&c;
		d(5) := input(12);
		d(4) := input(11);
		d(3) := input(10);
		d(2) := input(9);
		d(1) := input(8);
		d(0) := input(7);
		for i in 7 downto 1 loop
			if d(5) = '0' then
				for j in 4 downto 0 loop
				c(j) := d(j) xor '0';
				end loop;
			else
				for j in 4 downto 0 loop
				c(j) := d(j) xor p(j);
				end loop;
			end if;
			d := c&input(i-1);
		end loop;
		if d(5) = '0' then
				for j in 4 downto 0 loop
				c(j) := d(j) xor '0';
				end loop;
			else
				for j in 4 downto 0 loop
				c(j) := d(j) xor p(j);
				end loop;
			end if;
		o <= c;
		b_out <= o;
	end process;
END BEHAVIOR;
