-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 184 04/29/2009 Service Pack 1 SJ Web Edition
-- Created on Mon Nov 04 15:23:01 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY usb_download IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        rxf : IN STD_LOGIC := '0';
        rd : OUT STD_LOGIC
    );
END usb_download;

ARCHITECTURE BEHAVIOR OF usb_download IS
    TYPE type_fstate IS (wait_rxf_low,set_rd_low,latch_data_from_host);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= wait_rxf_low;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,rxf)
    BEGIN
        rd <= '0';
        CASE fstate IS
            WHEN wait_rxf_low =>
                IF (NOT((rxf = '1'))) THEN
                    reg_fstate <= set_rd_low;
                ELSIF ((rxf = '1')) THEN
                    reg_fstate <= wait_rxf_low;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= wait_rxf_low;
                END IF;

                rd <= '1';
            WHEN set_rd_low =>
                reg_fstate <= latch_data_from_host;

                rd <= '0';
            WHEN latch_data_from_host =>
                reg_fstate <= wait_rxf_low;
            WHEN OTHERS => 
                rd <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
