library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity mux8_1 is
port(	CIN: in std_logic_vector(7 downto 0);
		sel: in integer range 7 downto 0;
		COUT: out std_logic	);
end mux8_1;

architecture behav of mux8_1 is
COMPONENT multi_sel is
	generic( n: integer := 4	);
	port(	CIN: in std_logic_vector(n-1 downto 0);
			SEL: in integer range n-1 downto 0;
			COUT: out std_logic	);
end COMPONENT;

begin
	inst: multi_sel
		generic map(n =>8)
		port map(CIN =>CIN, COUT=>COUT, sel=>sel);
end behav;